

module MQ3(
  input         Alcohol_ent,                        
  output        Alcohol_sal
  );          

assign Alcohol_sal=Alcohol_ent;
endmodule

